lpm_dff5_inst : lpm_dff5 PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		q	 => q_sig
	);
