lpm_constant2_inst : lpm_constant2 PORT MAP (
		result	 => result_sig
	);
