lpm_inv0_inst : lpm_inv0 PORT MAP (
		data	 => data_sig,
		result	 => result_sig
	);
