lpm_constant3_inst : lpm_constant3 PORT MAP (
		result	 => result_sig
	);
